library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity data_ram is
    Port ( iCLK : in  STD_LOGIC;
           iRST : in  STD_LOGIC;
           iA : in  STD_LOGIC_VECTOR (7 downto 0); -- was 5 bits because the memory had 32 places
           iD : in  STD_LOGIC_VECTOR (31 downto 0);
           iWE : in  STD_LOGIC;
           oQ : out  STD_LOGIC_VECTOR (31 downto 0));
end data_ram;

architecture Behavioral of data_ram is

    type tMEM is array(0 to 255) of std_logic_vector(31 downto 0);
    signal rMEM : tMEM;
	 signal sMEM : tMEM := (others => x"00000000");

begin

    process (iCLK, iRST) begin
        if (iRST = '1') then
            for i in 0 to 255 loop
                rMEM(i) <= sMEM(i); 
            end loop;
        elsif (iCLK'event and iCLK = '1') then
            if (iWE = '1') then
                rMEM(to_integer(unsigned(iA))) <= iD;
            end if;
        end if;
    end process;
-- from here ---------------------------------------------------------------
 -- .data
	sMEM(0) 	<= "00000000000000000000000000000000";  -- _vrm
	sMEM(1) 	<= "00000000000000000000000000000000"; 
	sMEM(2) 	<= "00000000000000000000000000000000"; 
	sMEM(3) 	<= "00000000000000000000000000000000"; 
	sMEM(4) 	<= "00000000000000000000000000000000"; 
	sMEM(5) 	<= "00000000000000000000000000000000"; 
	sMEM(6) 	<= "00000000000000000000000000000000"; 
	sMEM(7) 	<= "00000000000000000000000000000000"; 
	sMEM(8) 	<= "00000000000000000000000000000000"; 
	sMEM(9) 	<= "00000000000000000000000000000000"; 
	sMEM(10) 	<= "00000000000000000000000000000000"; 
	sMEM(11) 	<= "00000000000000000000000000000000"; 
	sMEM(12) 	<= "00000000000000000000000000000000"; 
	sMEM(13) 	<= "00000000000000000000000000000000"; 
	sMEM(14) 	<= "00000000000000000000000000000000"; 
	sMEM(15) 	<= "00000000000000000000000000000000"; 
	sMEM(16) 	<= "00000000000000000000000000000000"; 
	sMEM(17) 	<= "00000000000000000000000000000000"; 
	sMEM(18) 	<= "00000000000000000000000000000000"; 
	sMEM(19) 	<= "00000000000000000000000000000000"; 
	sMEM(20) 	<= "00000000000000000000000000000000"; 
	sMEM(21) 	<= "00000000000000000000000000000000"; 
	sMEM(22) 	<= "00000000000000000000000000000000"; 
	sMEM(23) 	<= "00000000000000000000000000001111";  -- _m
	sMEM(24) 	<= "00000000000000000000000000000000";  -- _vtp
	sMEM(25) 	<= "00000000000000000000000000000000"; 
	sMEM(26) 	<= "00000000000000000000000000000000"; 
	sMEM(27) 	<= "00000000000000000000000000000000"; 
	sMEM(28) 	<= "00000000000000000000000000000000"; 
	sMEM(29) 	<= "00000000000000000000000000000000"; 
	sMEM(30) 	<= "00000000000000000000000000000000"; 
	sMEM(31) 	<= "00000000000000000000000000000000"; 
	sMEM(32) 	<= "00000000000000000000000000000000"; 
	sMEM(33) 	<= "00000000000000000000000000000000"; 
	sMEM(34) 	<= "00000000000000000000000000000000"; 
	sMEM(35) 	<= "00000000000000000000000000000000"; 
	sMEM(36) 	<= "11111111111111111111111111111101";  -- _t
--- to here  ---------------------------------------------------------------
    
oQ <= rMEM(to_integer(unsigned(iA)));

end Behavioral;
